`timescale 1ns / 1ps

module rModule_leds(
    input clk,
    input rst,
    output [1:0] led 
    );

endmodule
