`timescale 1ns / 1ps

module rModule_leds_2(
    input clk,
    input reset,
    input en,
    output [3:0] led
    );

endmodule